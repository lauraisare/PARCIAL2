library verilog;
use verilog.vl_types.all;
entity moore_peaje_vlg_vec_tst is
end moore_peaje_vlg_vec_tst;
