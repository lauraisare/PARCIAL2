library verilog;
use verilog.vl_types.all;
entity control_semaforo_vlg_vec_tst is
end control_semaforo_vlg_vec_tst;
