library verilog;
use verilog.vl_types.all;
entity categoria_vlg_vec_tst is
end categoria_vlg_vec_tst;
